module twiddle(
    input        [5:0]  idx,
    output logic [15:0] tw_re, // (16, 14)
    output logic [15:0] tw_im  // (16, 14)
);

logic [15:0] w_re[0:63];
logic [15:0] w_im[0:63];

/*
always_ff @(posedge clk) begin
    if (reset) begin
        tw_re <= #1 16'b0;
        tw_im <= #1 16'b0;
    end else begin
        tw_re <= #1 w_re[idx];
        tw_im <= #1 w_im[idx];
    end
end
*/

assign tw_re = w_re[idx];
assign tw_im = w_im[idx];

// cosine for real, sine for imag
assign w_re[0] = 16'b0100000000000000;		assign w_im[0] = 16'b0000000000000000;
assign w_re[1] = 16'b0011111110110001;		assign w_im[1] = 16'b1111100110111010;
assign w_re[2] = 16'b0011111011000101;		assign w_im[2] = 16'b1111001110000100;
assign w_re[3] = 16'b0011110100111111;		assign w_im[3] = 16'b1110110101101100;
assign w_re[4] = 16'b0011101100100001;		assign w_im[4] = 16'b1110011110000010;
assign w_re[5] = 16'b0011100001110001;		assign w_im[5] = 16'b1110000111010101;
assign w_re[6] = 16'b0011010100110111;		assign w_im[6] = 16'b1101110001110010;
assign w_re[7] = 16'b0011000101111001;		assign w_im[7] = 16'b1101011101100110;
assign w_re[8] = 16'b0010110101000001;		assign w_im[8] = 16'b1101001010111111;
assign w_re[9] = 16'b0010100010011010;		assign w_im[9] = 16'b1100111010000111;
assign w_re[10] = 16'b0010001110001110;		assign w_im[10] = 16'b1100101011001001;
assign w_re[11] = 16'b0001111000101011;		assign w_im[11] = 16'b1100011110001111;
assign w_re[12] = 16'b0001100001111110;		assign w_im[12] = 16'b1100010011011111;
assign w_re[13] = 16'b0001001010010100;		assign w_im[13] = 16'b1100001011000001;
assign w_re[14] = 16'b0000110001111100;		assign w_im[14] = 16'b1100000100111011;
assign w_re[15] = 16'b0000011001000110;		assign w_im[15] = 16'b1100000001001111;
assign w_re[16] = 16'b0000000000000000;		assign w_im[16] = 16'b1100000000000000;
assign w_re[17] = 16'b1111100110111010;		assign w_im[17] = 16'b1100000001001111;
assign w_re[18] = 16'b1111001110000100;		assign w_im[18] = 16'b1100000100111011;
assign w_re[19] = 16'b1110110101101100;		assign w_im[19] = 16'b1100001011000001;
assign w_re[20] = 16'b1110011110000010;		assign w_im[20] = 16'b1100010011011111;
assign w_re[21] = 16'b1110000111010101;		assign w_im[21] = 16'b1100011110001111;
assign w_re[22] = 16'b1101110001110010;		assign w_im[22] = 16'b1100101011001001;
assign w_re[23] = 16'b1101011101100110;		assign w_im[23] = 16'b1100111010000111;
assign w_re[24] = 16'b1101001010111111;		assign w_im[24] = 16'b1101001010111111;
assign w_re[25] = 16'b1100111010000111;		assign w_im[25] = 16'b1101011101100110;
assign w_re[26] = 16'b1100101011001001;		assign w_im[26] = 16'b1101110001110010;
assign w_re[27] = 16'b1100011110001111;		assign w_im[27] = 16'b1110000111010101;
assign w_re[28] = 16'b1100010011011111;		assign w_im[28] = 16'b1110011110000010;
assign w_re[29] = 16'b1100001011000001;		assign w_im[29] = 16'b1110110101101100;
assign w_re[30] = 16'b1100000100111011;		assign w_im[30] = 16'b1111001110000100;
assign w_re[31] = 16'b1100000001001111;		assign w_im[31] = 16'b1111100110111010;
assign w_re[32] = 16'b1100000000000000;		assign w_im[32] = 16'b0000000000000000;
assign w_re[33] = 16'b1100000001001111;		assign w_im[33] = 16'b0000011001000110;
assign w_re[34] = 16'b1100000100111011;		assign w_im[34] = 16'b0000110001111100;
assign w_re[35] = 16'b1100001011000001;		assign w_im[35] = 16'b0001001010010100;
assign w_re[36] = 16'b1100010011011111;		assign w_im[36] = 16'b0001100001111110;
assign w_re[37] = 16'b1100011110001111;		assign w_im[37] = 16'b0001111000101011;
assign w_re[38] = 16'b1100101011001001;		assign w_im[38] = 16'b0010001110001110;
assign w_re[39] = 16'b1100111010000111;		assign w_im[39] = 16'b0010100010011010;
assign w_re[40] = 16'b1101001010111111;		assign w_im[40] = 16'b0010110101000001;
assign w_re[41] = 16'b1101011101100110;		assign w_im[41] = 16'b0011000101111001;
assign w_re[42] = 16'b1101110001110010;		assign w_im[42] = 16'b0011010100110111;
assign w_re[43] = 16'b1110000111010101;		assign w_im[43] = 16'b0011100001110001;
assign w_re[44] = 16'b1110011110000010;		assign w_im[44] = 16'b0011101100100001;
assign w_re[45] = 16'b1110110101101100;		assign w_im[45] = 16'b0011110100111111;
assign w_re[46] = 16'b1111001110000100;		assign w_im[46] = 16'b0011111011000101;
assign w_re[47] = 16'b1111100110111010;		assign w_im[47] = 16'b0011111110110001;
assign w_re[48] = 16'b0000000000000000;		assign w_im[48] = 16'b0100000000000000;
assign w_re[49] = 16'b0000011001000110;		assign w_im[49] = 16'b0011111110110001;
assign w_re[50] = 16'b0000110001111100;		assign w_im[50] = 16'b0011111011000101;
assign w_re[51] = 16'b0001001010010100;		assign w_im[51] = 16'b0011110100111111;
assign w_re[52] = 16'b0001100001111110;		assign w_im[52] = 16'b0011101100100001;
assign w_re[53] = 16'b0001111000101011;		assign w_im[53] = 16'b0011100001110001;
assign w_re[54] = 16'b0010001110001110;		assign w_im[54] = 16'b0011010100110111;
assign w_re[55] = 16'b0010100010011010;		assign w_im[55] = 16'b0011000101111001;
assign w_re[56] = 16'b0010110101000001;		assign w_im[56] = 16'b0010110101000001;
assign w_re[57] = 16'b0011000101111001;		assign w_im[57] = 16'b0010100010011010;
assign w_re[58] = 16'b0011010100110111;		assign w_im[58] = 16'b0010001110001110;
assign w_re[59] = 16'b0011100001110001;		assign w_im[59] = 16'b0001111000101011;
assign w_re[60] = 16'b0011101100100001;		assign w_im[60] = 16'b0001100001111110;
assign w_re[61] = 16'b0011110100111111;		assign w_im[61] = 16'b0001001010010100;
assign w_re[62] = 16'b0011111011000101;		assign w_im[62] = 16'b0000110001111100;
assign w_re[63] = 16'b0011111110110001;		assign w_im[63] = 16'b0000011001000110;



endmodule
