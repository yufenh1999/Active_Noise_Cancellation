module hanning(
	input 		   clk,
	input 		   reset,
	input 		   in_valid,
	input 	signed [31:0] in_data, // fixed_point: (32,24)

	output	logic    	 out_valid,
	output 	logic signed [31:0] out_data 
);

	logic [6:0]  cnt, cnt_n;
	logic signed [63:0] temp;
	logic signed [31:0] LUT [63:0]; // fixed_point: (32,24)
	logic signed [31:0] out_data_n;

	assign LUT[0] = 32'b00000000000000000000000000000000;
	assign LUT[1] = 32'b00000000000000001010001011010100;
	assign LUT[2] = 32'b00000000000000101000100110110101;
	assign LUT[3] = 32'b00000000000001011010111111001010;
	assign LUT[4] = 32'b00000000000010100000110100010001;
	assign LUT[5] = 32'b00000000000011111001011001101111;
	assign LUT[6] = 32'b00000000000101100011110111001110;
	assign LUT[7] = 32'b00000000000111011111001001000001;
	assign LUT[8] = 32'b00000000001001101010000000101101;
	assign LUT[9] = 32'b00000000001100000011000101111100;
	assign LUT[10] = 32'b00000000001110101000110111011000;
	assign LUT[11] = 32'b00000000010001011001101011100011;
	assign LUT[12] = 32'b00000000010100010011110010000001;
	assign LUT[13] = 32'b00000000010111010101010100011001;
	assign LUT[14] = 32'b00000000011010011100010111100101;
	assign LUT[15] = 32'b00000000011101100110111100111110;
	assign LUT[16] = 32'b00000000100000110011000011101101;
	assign LUT[17] = 32'b00000000100011111110101001111110;
	assign LUT[18] = 32'b00000000100111000111101110010000;
	assign LUT[19] = 32'b00000000101010001100010000101011;
	assign LUT[20] = 32'b00000000101101001010010100001110;
	assign LUT[21] = 32'b00000000101111111111111111111111;
	assign LUT[22] = 32'b00000000110010101011100000011100;
	assign LUT[23] = 32'b00000000110101001011001000011111;
	assign LUT[24] = 32'b00000000110111011101010010100100;
	assign LUT[25] = 32'b00000000111001100000100001110000;
	assign LUT[26] = 32'b00000000111011010011100010100010;
	assign LUT[27] = 32'b00000000111100110101001011110010;
	assign LUT[28] = 32'b00000000111110000100011111011001;
	assign LUT[29] = 32'b00000000111111000000101010111001;
	assign LUT[30] = 32'b00000000111111101001001000000010;
	assign LUT[31] = 32'b00000000111111111101011101000100;
	assign LUT[32] = 32'b00000000111111111101011101000100;
	assign LUT[33] = 32'b00000000111111101001001000000010;
	assign LUT[34] = 32'b00000000111111000000101010111001;
	assign LUT[35] = 32'b00000000111110000100011111011001;
	assign LUT[36] = 32'b00000000111100110101001011110010;
	assign LUT[37] = 32'b00000000111011010011100010100010;
	assign LUT[38] = 32'b00000000111001100000100001110000;
	assign LUT[39] = 32'b00000000110111011101010010100100;
	assign LUT[40] = 32'b00000000110101001011001000011111;
	assign LUT[41] = 32'b00000000110010101011100000011100;
	assign LUT[42] = 32'b00000000101111111111111111111111;
	assign LUT[43] = 32'b00000000101101001010010100001110;
	assign LUT[44] = 32'b00000000101010001100010000101011;
	assign LUT[45] = 32'b00000000100111000111101110010000;
	assign LUT[46] = 32'b00000000100011111110101001111110;
	assign LUT[47] = 32'b00000000100000110011000011101101;
	assign LUT[48] = 32'b00000000011101100110111100111110;
	assign LUT[49] = 32'b00000000011010011100010111100101;
	assign LUT[50] = 32'b00000000010111010101010100011001;
	assign LUT[51] = 32'b00000000010100010011110010000001;
	assign LUT[52] = 32'b00000000010001011001101011100011;
	assign LUT[53] = 32'b00000000001110101000110111011000;
	assign LUT[54] = 32'b00000000001100000011000101111100;
	assign LUT[55] = 32'b00000000001001101010000000101101;
	assign LUT[56] = 32'b00000000000111011111001001000001;
	assign LUT[57] = 32'b00000000000101100011110111001110;
	assign LUT[58] = 32'b00000000000011111001011001101111;
	assign LUT[59] = 32'b00000000000010100000110100010001;
	assign LUT[60] = 32'b00000000000001011010111111001010;
	assign LUT[61] = 32'b00000000000000101000100110110101;
	assign LUT[62] = 32'b00000000000000001010001011010100;
	assign LUT[63] = 32'b00000000000000000000000000000000;




	always_comb begin
		cnt_n = cnt;
		if(in_valid) begin
			if(cnt == 7'd63) cnt_n = 0;
			else cnt_n = cnt + 1;
		end

		if(in_valid) temp = in_data * LUT[cnt];
		else temp = 0;

		out_data_n = temp[55:24];
		
	end

	always_ff @(posedge clk) begin
		if(reset) begin
			cnt <= 0;
			out_valid <= 0;
			out_data <= 0;
		end 
		else begin
			cnt <= cnt_n;
			out_valid <= in_valid;
			out_data <= out_data_n;
			
		end
	end 

endmodule
